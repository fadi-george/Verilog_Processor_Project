`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
//	Compare if two values are equal or not
//	
//////////////////////////////////////////////////////////////////////////////////
module Compar #(parameter M = 32) ( input [M-1:0] A , B,
												 output EqualD);

assign EqualD = (A == B) ? 1'b1 : 1'b0;		

endmodule
